package axil_pkg;
    typedef enum bit [1:0] {STATUS, CFG, TX, RX} register_t;
    typedef enum bit {WRITE, READ} rw_t;
endpackage: axil_pkg
